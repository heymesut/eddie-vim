// +FHDR----------------------------------------------------------------------------
// Project Name  : IC_Design
// Device        : Xilinx
// Author        : HonkW
// Email         : contact@honk.wang
// Website       : honk.wang
// Created On    : 2022/04/12 21:25
// Last Modified : 2022/04/12 21:25
// File Name     : test.v
// Description   :
//
// Copyright (c) 2022 NB Co.,Ltd..
// ALL RIGHTS RESERVED
//
// ---------------------------------------------------------------------------------
// Modification History:
// Date         By              Version                 Change Description
// ---------------------------------------------------------------------------------
// 2022/04/12   HonkW           1.0                     Original
// -FHDR----------------------------------------------------------------------------
`timescale 1ns/1ps

module test
(
clk
rst
);

endmodule

